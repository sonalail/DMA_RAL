`include "dma_intf.sv"
`include "ral_reg_block.sv"
`include "dma_seq_item.sv"
`include "dma_adapter.sv"
`include "dma_sequence.sv"
`include "dma_sequencer.sv"
`include "dma_driver.sv"
`include "dma_monitor.sv"
`include "dma_agent.sv"
`include "dma_scoreboard.sv"
`include "dma_environment.sv"
`include "dma_test.sv"
